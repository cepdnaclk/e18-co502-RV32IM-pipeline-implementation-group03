module cpu (

);







endmodule