module cpu (

);


// Stage 1 - Instruction Fetch





endmodule